@Filename: C:\vsm-lv\Lena\data\Salz\SH28\SH28-Hys-a000-RT.VHD
@Measurement Controlfilename: C:\vsm-lv\Stephie\Recipes\Hys-a000-RT.VHC
@Calibration filename: c:\vsm-lv\Stephie\settings\default.cal
@Parameter Filec:\vsm-lv\Stephie\settings\default.cal
@Operator: Lena
@Samplename: SH28
@Date: Tuesday, July 08, 2014    (2014-07-08)
@Time: 09:02:58
@Test ID: test
@Apparatus: EZ7;  Leibniz : MicroSense; first started on: Wednesday February 22, 2014
[Installed Options]
VSM Model="EZ7, EZ9 or EZ11"
VSM=TRUE    
Torque=FALSE    
Signal Processor="SR810"
Torque Signal Processor="NI-6210"
Unipolar=FALSE    
Automation=FALSE    
MR=FALSE    
Torque Signal Inversion=TRUE    
VSM DAQ Card=TRUE    
Time Constant="0.1 s"

[Signal and Coils]
Signal Connection="A-B"
Vector Coils=FALSE    
Stationary Coils=FALSE    
Z Coils=FALSE    
Sensor Angle="0 deg"
Time Between Averages=0.100000    
Y Averages Multiplier=1    
Reference Source="Internal"
SR830 Frequency=75.000000    

[Rotation]
Automatic Rotation=TRUE    
Rotate Option="Mdrive"
Rotation Display=FALSE    
Max Angle=400.000000    
Min Angle=-400.000000    
Rotation Serial Port=4    
Rotation Display Serial Port=1    
Torque Rotation Serial Port=4    

[Field]
Gaussmeter="FCM-10"
Gauss Probe="1 x"
Maximum Field=18000.000000    
Wait Time=0.000000    
Sweeprate Array="20.000, 50.000, 100.000, 200.000, 400.000, 500.000, 1000.000, 2000.000, 2000.000, 2000.000, "
Averaging Array="10, 5, 5, 2, 1, 1, 1, 1, 1, 1, "
Precision Array="0.010, 0.020, 0.050, 0.100, 0.100, 0.200, 0.200, 3.000, 3.000, 5.000, "
Stability Array="0.010, 0.020, 0.050, 0.100, 0.100, 0.200, 0.200, 3.000, 3.000, 5.000, "
FCM-10 Address="COM10"
Minimum Sweep Time=2.000000    
Minimum Sweep Rate Divider=100.000000    
Stability Time Between Readings=0.300000    
Number of Readings for Stability Check=4.000000    
Slow Approach=FALSE    
Slow Start %=100.000000    
Slow Approach Max Sweep Rate Divider=10.000000    
Max Slow Sweep Time=4.000000    

[MR]
MR Signal Processor=Manual VSM
Punch Through="Variable 0-10V"
Automation Comm Port=0
Max Current=20.000000    
Min AD Voltage=4.600000    
Max AD Voltage=7.000000    

[Temperature Control]
Temperature Control=TRUE    
Boil Off Nitrogen=FALSE    
Liquid Helium=FALSE    
Leave Temperature On=FALSE    
Temperature Control Type="SI 9700"
Sensor A="E-type"
Sensor B="E-type"
Control Sensor="A"
Sensor A Table=""
Sensor B Table=""
ITC Serial Port=2    
TC GPIB Address=15    
Temperature Log File="/c/vsm-lv/temperature.log"
Default Temperature=298.150000    
Gas Switching Temperature=333.150000    
Default Soak Time=120.000000    
Set Temperature Sample Time=10.000000    
Temperature Accuracy=1.000000    
Temperature Accuracy %=1.000000    
Automatic Gas Switching=FALSE    
1000 C Option=FALSE    
Number of points for accuracy wait=90    
Time between points for accuracy wait=1.000000    
Wait for Heat Exchanger Removal=FALSE    
Removal Temperature=0.000000    
Wait Time for Heat Exchanger Removal=0.000000    

[SI 9700]
P=1    
I=20    
D=0    
HE-P=1    
HE-I=20    
HE-D=0    
Max T Sweep Seed=1.000000
Min T Sweep Seed=0.200000
Max Heater Power=80    
Max T Sweep Speed=60.000000    
Min T Sweep Speed=12.000000    

[Other]
Transverse Direction="Absolute"
Default Transverse Direction=90.000000    
Time Dependence Start Field Distance=10.000000    
Minimum Remanence Wait Time=2.000000    
Default AC Demag Max Field=10000.000000    
AC Demag Minimum Field=1.000000    
Max Lockin Phase Error=90    
Mains Frequency=60.000000    
Samples Per Cycle=100    

[Interlock]
Door Lock=FALSE    
Interlock=FALSE    
Light Tower=FALSE    
Interlock Interface Name="Dev3"

[Torque Interface]
Torque Interface Name="Dev2"

[Exit Gas Heater Settings]
EGH PC Control=FALSE    
EGH Serial Port=0    
EGH Voltages=""

[VSM Interface]
VSM Interface Name="Dev1"

[MR Interface]
MR Interface Name="Dev1"

[DAQ Communication]
Protocol="Mx"
Remove Spikes=TRUE    

[Sensor Table]
1st Column=0    
Temperature Unit=0    

[Communication]
LIA 1 Address="COM5"
LIA 2 Address="COM5"
VSM Rotation Address="COM4"
Torque Rotation Address=""
Rotation Display Address=""
SI9700 Address="COM9"
EGH Address=""
Communication Mode="New"
LIA Baud Rate="19200"
LIA Serial Read Delay=50    

[LIA]
Local=0    
[FCM-10 Feedback Parameter Switching]
Switching = TRUE; Wait Before = 2000; Wait After = 1000; Progressive = TRUE; Progressive time =1.500000;
100 Oe: Field Setting Pars: FTCR = 10000; DR = 10000; DC = 10000; MDAC = 30000; Measurement Pars: FTCR = 100000; DR = 10000; DC = 10000; MDAC = 10000;
200 Oe: Field Setting Pars: FTCR = 5000; DR = 10000; DC = 10000; MDAC = 30000; Measurement Pars: FTCR = 50000; DR = 10000; DC = 10000; MDAC = 10000;
400 Oe: Field Setting Pars: FTCR = 5000; DR = 10000; DC = 10000; MDAC = 30000; Measurement Pars: FTCR = 50000; DR = 10000; DC = 10000; MDAC = 10000;
1k Oe: Field Setting Pars: FTCR = 5000; DR = 10000; DC = 10000; MDAC = 30000; Measurement Pars: FTCR = 50000; DR = 10000; DC = 10000; MDAC = 10000;
2 kOe: Field Setting Pars: FTCR = 5000; DR = 10000; DC = 10000; MDAC = 30000; Measurement Pars: FTCR = 20000; DR = 10000; DC = 10000; MDAC = 10000;
4 kOe: Field Setting Pars: FTCR = 1000; DR = 10000; DC = 10000; MDAC = 30000; Measurement Pars: FTCR = 20000; DR = 10000; DC = 10000; MDAC = 10000;
10 kOe: Field Setting Pars: FTCR = 500; DR = 10000; DC = 10000; MDAC = 30000; Measurement Pars: FTCR = 100000; DR = 10000; DC = 10000; MDAC = 10000;
20 kOe: Field Setting Pars: FTCR = 200; DR = 10000; DC = 1000; MDAC = 30000; Measurement Pars: FTCR = 100000; DR = 10000; DC = 1000; MDAC = 30000;
40 kOe: Field Setting Pars: FTCR = 100; DR = 10000; DC = 10000; MDAC = 30000; Measurement Pars: FTCR = 100000; DR = 10000; DC = 10000; MDAC = 30000;
100 kOe: Field Setting Pars: FTCR = 100; DR = 10000; DC = 10000; MDAC = 30000; Measurement Pars: FTCR = 100000; DR = 10000; DC = 10000; MDAC = 30000;
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 5.00 [mm] Volume : 1.963E-11 [m^3] Area = 1.963E+1 [mm^2] Mass = 2.722E-1 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: MicroSense EasyVSM Software version EasyVSM 20140521-01
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to -0.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Applied Field to -13999.7059 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Auto Range Signal to 13.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 7.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: -14000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 2000.0000 [Oe] Max Stepsize/Sweeprate = 2000.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Measured Signal(s) = X & Y
@Section 0 END
@Section 1: Hysteresis
@Preparation Actions: None
@Main Parameter Setup:
     From: -10000.0000 [Oe] To: -500.0000 [Oe] Min Stepsize/Sweeprate = 200.0000 [Oe] Max Stepsize/Sweeprate = 200.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: -500.0000 [Oe] To: 500.0000 [Oe] Min Stepsize/Sweeprate = 100.0000 [Oe] Max Stepsize/Sweeprate = 100.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: 500.0000 [Oe] To: 10000.0000 [Oe] Min Stepsize/Sweeprate = 200.0000 [Oe] Max Stepsize/Sweeprate = 200.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 18000.0000 [Oe] Min Stepsize/Sweeprate = 2000.0000 [Oe] Max Stepsize/Sweeprate = 2000.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 1
Plot 0: Hysteresis = On; Section: 0; Signal: X; Label: Hys X; Point style: 12; Interpolation: On; Color: 0; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = FALSE
Sensor Angle = 0 deg
@Gauss Range: 20 kOe
@Emu Range: 50 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 30
@Rot 0 deg cal: -21000
@Rot 360 deg cal: 21000
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 57.068
@Y Coils Correction Factor: 1.300
@Sample Shape Correction Factor: 1.000
@Coil Angle Alpha: 45.000
@Coil Angle Beta: -45.000
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 13
14999.670420   1.000000
15249.406962   1.000333
15500.452524   1.000604
15749.187630   1.000998
16000.025751   1.001472
16249.325953   1.001937
16500.206993   1.002473
16749.821932   1.002948
16999.837446   1.003547
17249.817193   1.004288
17499.847013   1.004968
17749.948363   1.005701
17999.527537   1.006649
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 0.000000
Background Subtraction = Yes   Method = Straight Line
Background slope x, y, z [emu/Oe] = -7.238824E-8   -0.000000E+0   0.000000E+0
Background Offset x, y, z [emu] = -2.131881E-6   -0.000000E+0   0.000000E+0
Angular Sensitivity Correction = Yes
Angular Sensitivity array length = 361
0.000000   1.000000E+0   0.000000E+0   0.000000
1.000000   9.999717E-1   0.000000E+0   0.000000
2.000000   9.999434E-1   0.000000E+0   0.000000
3.000000   9.999151E-1   0.000000E+0   0.000000
4.000000   9.998870E-1   0.000000E+0   0.000000
5.000000   9.998590E-1   0.000000E+0   0.000000
6.000000   9.998311E-1   0.000000E+0   0.000000
7.000000   9.998034E-1   0.000000E+0   0.000000
8.000000   9.997760E-1   0.000000E+0   0.000000
9.000000   9.997488E-1   0.000000E+0   0.000000
10.000000   9.997218E-1   0.000000E+0   0.000000
11.000000   9.996952E-1   0.000000E+0   0.000000
12.000000   9.996690E-1   0.000000E+0   0.000000
13.000000   9.996431E-1   0.000000E+0   0.000000
14.000000   9.996176E-1   0.000000E+0   0.000000
15.000000   9.995925E-1   0.000000E+0   0.000000
16.000000   9.995680E-1   0.000000E+0   0.000000
17.000000   9.995445E-1   0.000000E+0   0.000000
18.000000   9.995225E-1   0.000000E+0   0.000000
19.000000   9.995025E-1   0.000000E+0   0.000000
20.000000   9.994850E-1   0.000000E+0   0.000000
21.000000   9.994707E-1   0.000000E+0   0.000000
22.000000   9.994598E-1   0.000000E+0   0.000000
23.000000   9.994531E-1   0.000000E+0   0.000000
24.000000   9.994511E-1   0.000000E+0   0.000000
25.000000   9.994541E-1   0.000000E+0   0.000000
26.000000   9.994628E-1   0.000000E+0   0.000000
27.000000   9.994777E-1   0.000000E+0   0.000000
28.000000   9.994992E-1   0.000000E+0   0.000000
29.000000   9.995280E-1   0.000000E+0   0.000000
30.000000   9.995645E-1   0.000000E+0   0.000000
31.000000   9.996091E-1   0.000000E+0   0.000000
32.000000   9.996614E-1   0.000000E+0   0.000000
33.000000   9.997209E-1   0.000000E+0   0.000000
34.000000   9.997871E-1   0.000000E+0   0.000000
35.000000   9.998594E-1   0.000000E+0   0.000000
36.000000   9.999374E-1   0.000000E+0   0.000000
37.000000   1.000020E+0   0.000000E+0   0.000000
38.000000   1.000108E+0   0.000000E+0   0.000000
39.000000   1.000200E+0   0.000000E+0   0.000000
40.000000   1.000295E+0   0.000000E+0   0.000000
41.000000   1.000393E+0   0.000000E+0   0.000000
42.000000   1.000494E+0   0.000000E+0   0.000000
43.000000   1.000596E+0   0.000000E+0   0.000000
44.000000   1.000701E+0   0.000000E+0   0.000000
45.000000   1.000805E+0   0.000000E+0   0.000000
46.000000   1.000911E+0   0.000000E+0   0.000000
47.000000   1.001016E+0   0.000000E+0   0.000000
48.000000   1.001121E+0   0.000000E+0   0.000000
49.000000   1.001224E+0   0.000000E+0   0.000000
50.000000   1.001327E+0   0.000000E+0   0.000000
51.000000   1.001427E+0   0.000000E+0   0.000000
52.000000   1.001525E+0   0.000000E+0   0.000000
53.000000   1.001620E+0   0.000000E+0   0.000000
54.000000   1.001712E+0   0.000000E+0   0.000000
55.000000   1.001800E+0   0.000000E+0   0.000000
56.000000   1.001884E+0   0.000000E+0   0.000000
57.000000   1.001963E+0   0.000000E+0   0.000000
58.000000   1.002037E+0   0.000000E+0   0.000000
59.000000   1.002105E+0   0.000000E+0   0.000000
60.000000   1.002167E+0   0.000000E+0   0.000000
61.000000   1.002223E+0   0.000000E+0   0.000000
62.000000   1.002273E+0   0.000000E+0   0.000000
63.000000   1.002317E+0   0.000000E+0   0.000000
64.000000   1.002357E+0   0.000000E+0   0.000000
65.000000   1.002392E+0   0.000000E+0   0.000000
66.000000   1.002423E+0   0.000000E+0   0.000000
67.000000   1.002451E+0   0.000000E+0   0.000000
68.000000   1.002476E+0   0.000000E+0   0.000000
69.000000   1.002498E+0   0.000000E+0   0.000000
70.000000   1.002519E+0   0.000000E+0   0.000000
71.000000   1.002538E+0   0.000000E+0   0.000000
72.000000   1.002557E+0   0.000000E+0   0.000000
73.000000   1.002575E+0   0.000000E+0   0.000000
74.000000   1.002594E+0   0.000000E+0   0.000000
75.000000   1.002614E+0   0.000000E+0   0.000000
76.000000   1.002634E+0   0.000000E+0   0.000000
77.000000   1.002656E+0   0.000000E+0   0.000000
78.000000   1.002678E+0   0.000000E+0   0.000000
79.000000   1.002700E+0   0.000000E+0   0.000000
80.000000   1.002722E+0   0.000000E+0   0.000000
81.000000   1.002742E+0   0.000000E+0   0.000000
82.000000   1.002762E+0   0.000000E+0   0.000000
83.000000   1.002779E+0   0.000000E+0   0.000000
84.000000   1.002795E+0   0.000000E+0   0.000000
85.000000   1.002808E+0   0.000000E+0   0.000000
86.000000   1.002817E+0   0.000000E+0   0.000000
87.000000   1.002823E+0   0.000000E+0   0.000000
88.000000   1.002825E+0   0.000000E+0   0.000000
89.000000   1.002823E+0   0.000000E+0   0.000000
90.000000   1.002816E+0   0.000000E+0   0.000000
91.000000   1.002803E+0   0.000000E+0   0.000000
92.000000   1.002783E+0   0.000000E+0   0.000000
93.000000   1.002752E+0   0.000000E+0   0.000000
94.000000   1.002709E+0   0.000000E+0   0.000000
95.000000   1.002651E+0   0.000000E+0   0.000000
96.000000   1.002576E+0   0.000000E+0   0.000000
97.000000   1.002482E+0   0.000000E+0   0.000000
98.000000   1.002365E+0   0.000000E+0   0.000000
99.000000   1.002224E+0   0.000000E+0   0.000000
100.000000   1.002057E+0   0.000000E+0   0.000000
101.000000   1.001860E+0   0.000000E+0   0.000000
102.000000   1.001632E+0   0.000000E+0   0.000000
103.000000   1.001370E+0   0.000000E+0   0.000000
104.000000   1.001072E+0   0.000000E+0   0.000000
105.000000   1.000735E+0   0.000000E+0   0.000000
106.000000   1.000359E+0   0.000000E+0   0.000000
107.000000   9.999441E-1   0.000000E+0   0.000000
108.000000   9.994949E-1   0.000000E+0   0.000000
109.000000   9.990141E-1   0.000000E+0   0.000000
110.000000   9.985049E-1   0.000000E+0   0.000000
111.000000   9.979705E-1   0.000000E+0   0.000000
112.000000   9.974140E-1   0.000000E+0   0.000000
113.000000   9.968386E-1   0.000000E+0   0.000000
114.000000   9.962473E-1   0.000000E+0   0.000000
115.000000   9.956433E-1   0.000000E+0   0.000000
116.000000   9.950298E-1   0.000000E+0   0.000000
117.000000   9.944099E-1   0.000000E+0   0.000000
118.000000   9.937868E-1   0.000000E+0   0.000000
119.000000   9.931635E-1   0.000000E+0   0.000000
120.000000   9.925432E-1   0.000000E+0   0.000000
121.000000   9.919287E-1   0.000000E+0   0.000000
122.000000   9.913204E-1   0.000000E+0   0.000000
123.000000   9.907185E-1   0.000000E+0   0.000000
124.000000   9.901232E-1   0.000000E+0   0.000000
125.000000   9.895345E-1   0.000000E+0   0.000000
126.000000   9.889526E-1   0.000000E+0   0.000000
127.000000   9.883776E-1   0.000000E+0   0.000000
128.000000   9.878096E-1   0.000000E+0   0.000000
129.000000   9.872488E-1   0.000000E+0   0.000000
130.000000   9.866951E-1   0.000000E+0   0.000000
131.000000   9.861489E-1   0.000000E+0   0.000000
132.000000   9.856102E-1   0.000000E+0   0.000000
133.000000   9.850790E-1   0.000000E+0   0.000000
134.000000   9.845556E-1   0.000000E+0   0.000000
135.000000   9.840401E-1   0.000000E+0   0.000000
136.000000   9.835323E-1   0.000000E+0   0.000000
137.000000   9.830315E-1   0.000000E+0   0.000000
138.000000   9.825365E-1   0.000000E+0   0.000000
139.000000   9.820462E-1   0.000000E+0   0.000000
140.000000   9.815598E-1   0.000000E+0   0.000000
141.000000   9.810760E-1   0.000000E+0   0.000000
142.000000   9.805938E-1   0.000000E+0   0.000000
143.000000   9.801121E-1   0.000000E+0   0.000000
144.000000   9.796299E-1   0.000000E+0   0.000000
145.000000   9.791462E-1   0.000000E+0   0.000000
146.000000   9.786598E-1   0.000000E+0   0.000000
147.000000   9.781697E-1   0.000000E+0   0.000000
148.000000   9.776749E-1   0.000000E+0   0.000000
149.000000   9.771742E-1   0.000000E+0   0.000000
150.000000   9.766667E-1   0.000000E+0   0.000000
151.000000   9.761516E-1   0.000000E+0   0.000000
152.000000   9.756301E-1   0.000000E+0   0.000000
153.000000   9.751034E-1   0.000000E+0   0.000000
154.000000   9.745730E-1   0.000000E+0   0.000000
155.000000   9.740404E-1   0.000000E+0   0.000000
156.000000   9.735069E-1   0.000000E+0   0.000000
157.000000   9.729740E-1   0.000000E+0   0.000000
158.000000   9.724431E-1   0.000000E+0   0.000000
159.000000   9.719156E-1   0.000000E+0   0.000000
160.000000   9.713929E-1   0.000000E+0   0.000000
161.000000   9.708765E-1   0.000000E+0   0.000000
162.000000   9.703678E-1   0.000000E+0   0.000000
163.000000   9.698681E-1   0.000000E+0   0.000000
164.000000   9.693790E-1   0.000000E+0   0.000000
165.000000   9.689018E-1   0.000000E+0   0.000000
166.000000   9.684377E-1   0.000000E+0   0.000000
167.000000   9.679871E-1   0.000000E+0   0.000000
168.000000   9.675501E-1   0.000000E+0   0.000000
169.000000   9.671268E-1   0.000000E+0   0.000000
170.000000   9.667174E-1   0.000000E+0   0.000000
171.000000   9.663220E-1   0.000000E+0   0.000000
172.000000   9.659408E-1   0.000000E+0   0.000000
173.000000   9.655737E-1   0.000000E+0   0.000000
174.000000   9.652211E-1   0.000000E+0   0.000000
175.000000   9.648829E-1   0.000000E+0   0.000000
176.000000   9.645594E-1   0.000000E+0   0.000000
177.000000   9.642507E-1   0.000000E+0   0.000000
178.000000   9.639568E-1   0.000000E+0   0.000000
179.000000   9.636780E-1   0.000000E+0   0.000000
180.000000   9.634143E-1   0.000000E+0   0.000000
181.000000   9.631659E-1   0.000000E+0   0.000000
182.000000   9.629324E-1   0.000000E+0   0.000000
183.000000   9.627136E-1   0.000000E+0   0.000000
184.000000   9.625093E-1   0.000000E+0   0.000000
185.000000   9.623191E-1   0.000000E+0   0.000000
186.000000   9.621427E-1   0.000000E+0   0.000000
187.000000   9.619798E-1   0.000000E+0   0.000000
188.000000   9.618302E-1   0.000000E+0   0.000000
189.000000   9.616936E-1   0.000000E+0   0.000000
190.000000   9.615697E-1   0.000000E+0   0.000000
191.000000   9.614581E-1   0.000000E+0   0.000000
192.000000   9.613587E-1   0.000000E+0   0.000000
193.000000   9.612710E-1   0.000000E+0   0.000000
194.000000   9.611949E-1   0.000000E+0   0.000000
195.000000   9.611300E-1   0.000000E+0   0.000000
196.000000   9.610762E-1   0.000000E+0   0.000000
197.000000   9.610335E-1   0.000000E+0   0.000000
198.000000   9.610023E-1   0.000000E+0   0.000000
199.000000   9.609828E-1   0.000000E+0   0.000000
200.000000   9.609752E-1   0.000000E+0   0.000000
201.000000   9.609798E-1   0.000000E+0   0.000000
202.000000   9.609968E-1   0.000000E+0   0.000000
203.000000   9.610265E-1   0.000000E+0   0.000000
204.000000   9.610691E-1   0.000000E+0   0.000000
205.000000   9.611249E-1   0.000000E+0   0.000000
206.000000   9.611942E-1   0.000000E+0   0.000000
207.000000   9.612771E-1   0.000000E+0   0.000000
208.000000   9.613739E-1   0.000000E+0   0.000000
209.000000   9.614849E-1   0.000000E+0   0.000000
210.000000   9.616103E-1   0.000000E+0   0.000000
211.000000   9.617504E-1   0.000000E+0   0.000000
212.000000   9.619054E-1   0.000000E+0   0.000000
213.000000   9.620756E-1   0.000000E+0   0.000000
214.000000   9.622612E-1   0.000000E+0   0.000000
215.000000   9.624626E-1   0.000000E+0   0.000000
216.000000   9.626800E-1   0.000000E+0   0.000000
217.000000   9.629136E-1   0.000000E+0   0.000000
218.000000   9.631637E-1   0.000000E+0   0.000000
219.000000   9.634307E-1   0.000000E+0   0.000000
220.000000   9.637146E-1   0.000000E+0   0.000000
221.000000   9.640159E-1   0.000000E+0   0.000000
222.000000   9.643348E-1   0.000000E+0   0.000000
223.000000   9.646715E-1   0.000000E+0   0.000000
224.000000   9.650264E-1   0.000000E+0   0.000000
225.000000   9.653996E-1   0.000000E+0   0.000000
226.000000   9.657914E-1   0.000000E+0   0.000000
227.000000   9.662019E-1   0.000000E+0   0.000000
228.000000   9.666311E-1   0.000000E+0   0.000000
229.000000   9.670791E-1   0.000000E+0   0.000000
230.000000   9.675458E-1   0.000000E+0   0.000000
231.000000   9.680314E-1   0.000000E+0   0.000000
232.000000   9.685358E-1   0.000000E+0   0.000000
233.000000   9.690591E-1   0.000000E+0   0.000000
234.000000   9.696013E-1   0.000000E+0   0.000000
235.000000   9.701625E-1   0.000000E+0   0.000000
236.000000   9.707427E-1   0.000000E+0   0.000000
237.000000   9.713419E-1   0.000000E+0   0.000000
238.000000   9.719602E-1   0.000000E+0   0.000000
239.000000   9.725976E-1   0.000000E+0   0.000000
240.000000   9.732541E-1   0.000000E+0   0.000000
241.000000   9.739297E-1   0.000000E+0   0.000000
242.000000   9.746244E-1   0.000000E+0   0.000000
243.000000   9.753379E-1   0.000000E+0   0.000000
244.000000   9.760701E-1   0.000000E+0   0.000000
245.000000   9.768209E-1   0.000000E+0   0.000000
246.000000   9.775899E-1   0.000000E+0   0.000000
247.000000   9.783772E-1   0.000000E+0   0.000000
248.000000   9.791825E-1   0.000000E+0   0.000000
249.000000   9.800057E-1   0.000000E+0   0.000000
250.000000   9.808465E-1   0.000000E+0   0.000000
251.000000   9.817049E-1   0.000000E+0   0.000000
252.000000   9.825807E-1   0.000000E+0   0.000000
253.000000   9.834737E-1   0.000000E+0   0.000000
254.000000   9.843837E-1   0.000000E+0   0.000000
255.000000   9.853107E-1   0.000000E+0   0.000000
256.000000   9.862538E-1   0.000000E+0   0.000000
257.000000   9.872100E-1   0.000000E+0   0.000000
258.000000   9.881759E-1   0.000000E+0   0.000000
259.000000   9.891479E-1   0.000000E+0   0.000000
260.000000   9.901225E-1   0.000000E+0   0.000000
261.000000   9.910960E-1   0.000000E+0   0.000000
262.000000   9.920650E-1   0.000000E+0   0.000000
263.000000   9.930260E-1   0.000000E+0   0.000000
264.000000   9.939753E-1   0.000000E+0   0.000000
265.000000   9.949095E-1   0.000000E+0   0.000000
266.000000   9.958250E-1   0.000000E+0   0.000000
267.000000   9.967182E-1   0.000000E+0   0.000000
268.000000   9.975857E-1   0.000000E+0   0.000000
269.000000   9.984238E-1   0.000000E+0   0.000000
270.000000   9.992290E-1   0.000000E+0   0.000000
271.000000   9.999985E-1   0.000000E+0   0.000000
272.000000   1.000732E+0   0.000000E+0   0.000000
273.000000   1.001430E+0   0.000000E+0   0.000000
274.000000   1.002093E+0   0.000000E+0   0.000000
275.000000   1.002722E+0   0.000000E+0   0.000000
276.000000   1.003316E+0   0.000000E+0   0.000000
277.000000   1.003877E+0   0.000000E+0   0.000000
278.000000   1.004405E+0   0.000000E+0   0.000000
279.000000   1.004900E+0   0.000000E+0   0.000000
280.000000   1.005363E+0   0.000000E+0   0.000000
281.000000   1.005794E+0   0.000000E+0   0.000000
282.000000   1.006194E+0   0.000000E+0   0.000000
283.000000   1.006563E+0   0.000000E+0   0.000000
284.000000   1.006902E+0   0.000000E+0   0.000000
285.000000   1.007211E+0   0.000000E+0   0.000000
286.000000   1.007491E+0   0.000000E+0   0.000000
287.000000   1.007743E+0   0.000000E+0   0.000000
288.000000   1.007968E+0   0.000000E+0   0.000000
289.000000   1.008168E+0   0.000000E+0   0.000000
290.000000   1.008345E+0   0.000000E+0   0.000000
291.000000   1.008499E+0   0.000000E+0   0.000000
292.000000   1.008632E+0   0.000000E+0   0.000000
293.000000   1.008747E+0   0.000000E+0   0.000000
294.000000   1.008843E+0   0.000000E+0   0.000000
295.000000   1.008922E+0   0.000000E+0   0.000000
296.000000   1.008987E+0   0.000000E+0   0.000000
297.000000   1.009038E+0   0.000000E+0   0.000000
298.000000   1.009076E+0   0.000000E+0   0.000000
299.000000   1.009104E+0   0.000000E+0   0.000000
300.000000   1.009123E+0   0.000000E+0   0.000000
301.000000   1.009133E+0   0.000000E+0   0.000000
302.000000   1.009136E+0   0.000000E+0   0.000000
303.000000   1.009133E+0   0.000000E+0   0.000000
304.000000   1.009124E+0   0.000000E+0   0.000000
305.000000   1.009110E+0   0.000000E+0   0.000000
306.000000   1.009093E+0   0.000000E+0   0.000000
307.000000   1.009072E+0   0.000000E+0   0.000000
308.000000   1.009048E+0   0.000000E+0   0.000000
309.000000   1.009023E+0   0.000000E+0   0.000000
310.000000   1.008996E+0   0.000000E+0   0.000000
311.000000   1.008970E+0   0.000000E+0   0.000000
312.000000   1.008944E+0   0.000000E+0   0.000000
313.000000   1.008919E+0   0.000000E+0   0.000000
314.000000   1.008896E+0   0.000000E+0   0.000000
315.000000   1.008877E+0   0.000000E+0   0.000000
316.000000   1.008861E+0   0.000000E+0   0.000000
317.000000   1.008848E+0   0.000000E+0   0.000000
318.000000   1.008838E+0   0.000000E+0   0.000000
319.000000   1.008830E+0   0.000000E+0   0.000000
320.000000   1.008824E+0   0.000000E+0   0.000000
321.000000   1.008820E+0   0.000000E+0   0.000000
322.000000   1.008817E+0   0.000000E+0   0.000000
323.000000   1.008815E+0   0.000000E+0   0.000000
324.000000   1.008813E+0   0.000000E+0   0.000000
325.000000   1.008810E+0   0.000000E+0   0.000000
326.000000   1.008808E+0   0.000000E+0   0.000000
327.000000   1.008804E+0   0.000000E+0   0.000000
328.000000   1.008799E+0   0.000000E+0   0.000000
329.000000   1.008792E+0   0.000000E+0   0.000000
330.000000   1.008782E+0   0.000000E+0   0.000000
331.000000   1.008770E+0   0.000000E+0   0.000000
332.000000   1.008755E+0   0.000000E+0   0.000000
333.000000   1.008735E+0   0.000000E+0   0.000000
334.000000   1.008709E+0   0.000000E+0   0.000000
335.000000   1.008677E+0   0.000000E+0   0.000000
336.000000   1.008638E+0   0.000000E+0   0.000000
337.000000   1.008590E+0   0.000000E+0   0.000000
338.000000   1.008533E+0   0.000000E+0   0.000000
339.000000   1.008467E+0   0.000000E+0   0.000000
340.000000   1.008389E+0   0.000000E+0   0.000000
341.000000   1.008299E+0   0.000000E+0   0.000000
342.000000   1.008196E+0   0.000000E+0   0.000000
343.000000   1.008080E+0   0.000000E+0   0.000000
344.000000   1.007949E+0   0.000000E+0   0.000000
345.000000   1.007802E+0   0.000000E+0   0.000000
346.000000   1.007640E+0   0.000000E+0   0.000000
347.000000   1.007461E+0   0.000000E+0   0.000000
348.000000   1.007269E+0   0.000000E+0   0.000000
349.000000   1.007063E+0   0.000000E+0   0.000000
350.000000   1.006845E+0   0.000000E+0   0.000000
351.000000   1.006616E+0   0.000000E+0   0.000000
352.000000   1.006377E+0   0.000000E+0   0.000000
353.000000   1.006129E+0   0.000000E+0   0.000000
354.000000   1.005873E+0   0.000000E+0   0.000000
355.000000   1.005611E+0   0.000000E+0   0.000000
356.000000   1.005343E+0   0.000000E+0   0.000000
357.000000   1.005071E+0   0.000000E+0   0.000000
358.000000   1.004796E+0   0.000000E+0   0.000000
359.000000   1.004518E+0   0.000000E+0   0.000000
360.000000   1.004240E+0   0.000000E+0   0.000000
Remove Slope = Yes    Slope Correction Start Field = 0.000 [Oe], Use Max Field = Yes, Slopealculation Max Field = 18000.000 [Oe]
Remove Signal Offset = No
Remove Signal Drift = FALSE; Drift # Points = 0
Remove Field Offset = No
Field Offset Method = Automatic
Field Offset = 0.0000
Remove Field Lag = No
Field Lag Method = Automatic
Field Lag = 0.0000
Cubic Spline Interpolation = No   # Points = 100
Noise Filter = No   Filter Order = 20   Filter Type = Median
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 1.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = Monday, July 07, 2014  09:20:29
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Temperature 2, Sample Temperature [degC]
Column 4: Raw Applied Field, Applied Field [Oe]
Column 5: Applied Field, Applied Field [Oe]
Column 6: Field Angle, Field Angle [deg]
Column 7: Raw Applied Field For Plot , Applied Field [Oe]
Column 8: Applied Field For Plot , Applied Field [Oe]
Column 9: Raw Signal Mx, Moment as measured [memu]
Column 10: Raw Signal My, Moment as measured [memu]
Column 11: Signal X direction, Moment [emu]
Column 12: Signal Y direction, Moment [emu]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Temperature_2   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction      
@Time at start of measurement: 09:02:59
@@Data
New Section: Section 0: 
1.453500E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.399982E+4   -1.399982E+4   -1.161182E+0   0.000000E+0   -2.172473E-3   0.000000E+0   
2.907600E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.199999E+4   -1.199999E+4   -1.106947E+0   0.000000E+0   -1.973473E-3   0.000000E+0   
4.646500E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.000024E+4   -1.000024E+4   -1.059563E+0   0.000000E+0   -1.781330E-3   0.000000E+0   
6.173500E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.800147E+3   -9.800147E+3   -1.048243E+0   0.000000E+0   -1.755526E-3   0.000000E+0   
7.372300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.600204E+3   -9.600204E+3   -1.039898E+0   0.000000E+0   -1.732708E-3   0.000000E+0   
8.566300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.400146E+3   -9.400146E+3   -1.034825E+0   0.000000E+0   -1.713153E-3   0.000000E+0   
9.759500E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.200167E+3   -9.200167E+3   -1.030623E+0   0.000000E+0   -1.694475E-3   0.000000E+0   
1.094890E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.000099E+3   -9.000099E+3   -1.024911E+0   0.000000E+0   -1.674280E-3   0.000000E+0   
1.213770E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.800020E+3   -8.800020E+3   -1.020124E+0   0.000000E+0   -1.655010E-3   0.000000E+0   
1.333700E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.600163E+3   -8.600163E+3   -1.014132E+0   0.000000E+0   -1.634551E-3   0.000000E+0   
1.453090E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.400180E+3   -8.400180E+3   -1.008934E+0   0.000000E+0   -1.614877E-3   0.000000E+0   
1.572460E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.200187E+3   -8.200187E+3   -1.000526E+0   0.000000E+0   -1.591991E-3   0.000000E+0   
1.691350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.000187E+3   -8.000187E+3   -9.954341E-1   0.000000E+0   -1.572422E-3   0.000000E+0   
1.810760E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.800201E+3   -7.800201E+3   -9.859596E-1   0.000000E+0   -1.548471E-3   0.000000E+0   
1.929640E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.600193E+3   -7.600193E+3   -9.827071E-1   0.000000E+0   -1.530740E-3   0.000000E+0   
2.049530E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.400190E+3   -7.400190E+3   -9.745225E-1   0.000000E+0   -1.508077E-3   0.000000E+0   
2.168960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.200254E+3   -7.200254E+3   -9.697457E-1   0.000000E+0   -1.488828E-3   0.000000E+0   
2.288350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.000128E+3   -7.000128E+3   -9.621676E-1   0.000000E+0   -1.466763E-3   0.000000E+0   
2.407780E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.800085E+3   -6.800085E+3   -9.558074E-1   0.000000E+0   -1.445922E-3   0.000000E+0   
2.527790E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.600138E+3   -6.600138E+3   -9.479659E-1   0.000000E+0   -1.423606E-3   0.000000E+0   
2.647310E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.400242E+3   -6.400242E+3   -9.418150E-1   0.000000E+0   -1.402985E-3   0.000000E+0   
2.766830E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.200156E+3   -6.200156E+3   -9.365604E-1   0.000000E+0   -1.383247E-3   0.000000E+0   
2.886350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.999998E+3   -5.999998E+3   -9.263450E-1   0.000000E+0   -1.358542E-3   0.000000E+0   
3.005840E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.800137E+3   -5.800137E+3   -9.211299E-1   0.000000E+0   -1.338860E-3   0.000000E+0   
3.125350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.600137E+3   -5.600137E+3   -9.105529E-1   0.000000E+0   -1.313805E-3   0.000000E+0   
3.244820E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.400026E+3   -5.400026E+3   -9.039486E-1   0.000000E+0   -1.292715E-3   0.000000E+0   
3.363850E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.200029E+3   -5.200029E+3   -8.969259E-1   0.000000E+0   -1.271215E-3   0.000000E+0   
3.483340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.000122E+3   -5.000122E+3   -8.889644E-1   0.000000E+0   -1.248783E-3   0.000000E+0   
3.602830E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.800043E+3   -4.800043E+3   -8.807722E-1   0.000000E+0   -1.226107E-3   0.000000E+0   
3.722340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.599999E+3   -4.599999E+3   -8.717974E-1   0.000000E+0   -1.202651E-3   0.000000E+0   
3.841340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.400078E+3   -4.400078E+3   -8.616852E-1   0.000000E+0   -1.178067E-3   0.000000E+0   
3.960860E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.199920E+3   -4.199920E+3   -8.523383E-1   0.000000E+0   -1.154231E-3   0.000000E+0   
4.080380E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.000027E+3   -4.000027E+3   -8.426935E-1   0.000000E+0   -1.130117E-3   0.000000E+0   
4.199910E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.800102E+3   -3.800102E+3   -8.317027E-1   0.000000E+0   -1.104654E-3   0.000000E+0   
4.319390E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.600044E+3   -3.600044E+3   -8.243541E-1   0.000000E+0   -1.082823E-3   0.000000E+0   
4.438910E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.399865E+3   -3.399865E+3   -8.096039E-1   0.000000E+0   -1.053582E-3   0.000000E+0   
4.558440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.200037E+3   -3.200037E+3   -7.974500E-1   0.000000E+0   -1.026963E-3   0.000000E+0   
4.677950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.000054E+3   -3.000054E+3   -7.852967E-1   0.000000E+0   -1.000334E-3   0.000000E+0   
4.797470E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.799954E+3   -2.799954E+3   -7.726228E-1   0.000000E+0   -9.731747E-4   0.000000E+0   
4.916970E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.600107E+3   -2.600107E+3   -7.603814E-1   0.000000E+0   -9.464668E-4   0.000000E+0   
5.036490E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.399867E+3   -2.399867E+3   -7.407769E-1   0.000000E+0   -9.123672E-4   0.000000E+0   
5.156000E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.199992E+3   -2.199992E+3   -7.228554E-1   0.000000E+0   -8.799771E-4   0.000000E+0   
5.276010E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.999931E+3   -1.999931E+3   -7.013866E-1   0.000000E+0   -8.440262E-4   0.000000E+0   
5.394020E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.799927E+3   -1.799927E+3   -6.802227E-1   0.000000E+0   -8.083844E-4   0.000000E+0   
5.513050E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.599884E+3   -1.599884E+3   -6.574467E-1   0.000000E+0   -7.711276E-4   0.000000E+0   
5.632050E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.400077E+3   -1.400077E+3   -6.274967E-1   0.000000E+0   -7.267139E-4   0.000000E+0   
5.751080E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.200030E+3   -1.200030E+3   -5.912459E-1   0.000000E+0   -6.759821E-4   0.000000E+0   
5.870090E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.998903E+2   -9.998903E+2   -5.564513E-1   0.000000E+0   -6.266997E-4   0.000000E+0   
5.988590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.999150E+2   -7.999150E+2   -5.104817E-1   0.000000E+0   -5.662543E-4   0.000000E+0   
6.107100E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.000578E+2   -6.000578E+2   -4.610431E-1   0.000000E+0   -5.023484E-4   0.000000E+0   
6.225100E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.998824E+2   -4.998824E+2   -4.297478E-1   0.000000E+0   -4.638015E-4   0.000000E+0   
6.375990E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.998894E+2   -3.998894E+2   -3.982557E-1   0.000000E+0   -4.250711E-4   0.000000E+0   
6.494010E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.998606E+2   -2.998606E+2   -3.632133E-1   0.000000E+0   -3.827878E-4   0.000000E+0   
6.612020E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.000107E+2   -2.000107E+2   -3.218639E-1   0.000000E+0   -3.342105E-4   0.000000E+0   
6.730040E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.992111E+1   -9.992111E+1   -2.736762E-1   0.000000E+0   -2.787774E-4   0.000000E+0   
6.848050E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.326898E-1   1.326898E-1   -2.119880E-1   0.000000E+0   -2.098465E-4   0.000000E+0   
6.971580E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.001579E+2   1.001579E+2   -1.397311E-1   0.000000E+0   -1.303490E-4   0.000000E+0   
7.095110E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.000328E+2   2.000328E+2   -7.114466E-2   0.000000E+0   -5.453276E-5   0.000000E+0   
7.215150E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.000866E+2   3.000866E+2   -7.578984E-3   0.000000E+0   1.627564E-5   0.000000E+0   
7.338690E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.001655E+2   4.001655E+2   5.051231E-2   0.000000E+0   8.161146E-5   0.000000E+0   
7.458710E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.002193E+2   5.002193E+2   9.919279E-2   0.000000E+0   1.375347E-4   0.000000E+0   
7.615590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.002196E+2   7.002196E+2   1.791317E-1   0.000000E+0   2.319512E-4   0.000000E+0   
7.740120E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.000303E+2   9.000303E+2   2.448167E-1   0.000000E+0   3.121002E-4   0.000000E+0   
7.864650E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.100016E+3   1.100016E+3   2.979153E-1   0.000000E+0   3.796754E-4   0.000000E+0   
7.989180E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.300149E+3   1.300149E+3   3.398032E-1   0.000000E+0   4.360506E-4   0.000000E+0   
8.113710E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.499967E+3   1.499967E+3   3.793526E-1   0.000000E+0   4.900644E-4   0.000000E+0   
8.238240E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.700071E+3   1.700071E+3   4.138671E-1   0.000000E+0   5.390641E-4   0.000000E+0   
8.362840E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.900271E+3   1.900271E+3   4.454105E-1   0.000000E+0   5.850997E-4   0.000000E+0   
8.488360E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.100136E+3   2.100136E+3   4.743196E-1   0.000000E+0   6.284766E-4   0.000000E+0   
8.614380E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.300057E+3   2.300057E+3   4.980307E-1   0.000000E+0   6.666597E-4   0.000000E+0   
8.739400E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.500076E+3   2.500076E+3   5.208845E-1   0.000000E+0   7.039925E-4   0.000000E+0   
8.864450E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.700147E+3   2.700147E+3   5.482594E-1   0.000000E+0   7.458502E-4   0.000000E+0   
8.989500E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.900234E+3   2.900234E+3   5.692744E-1   0.000000E+0   7.813491E-4   0.000000E+0   
9.114530E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.100137E+3   3.100137E+3   5.869866E-1   0.000000E+0   8.135320E-4   0.000000E+0   
9.239580E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.299991E+3   3.299991E+3   6.064780E-1   0.000000E+0   8.474904E-4   0.000000E+0   
9.364590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.500299E+3   3.500299E+3   6.251796E-1   0.000000E+0   8.806920E-4   0.000000E+0   
9.489590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.700224E+3   3.700224E+3   6.443134E-1   0.000000E+0   9.142980E-4   0.000000E+0   
9.614560E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.900114E+3   3.900114E+3   6.607739E-1   0.000000E+0   9.452282E-4   0.000000E+0   
9.740040E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.100225E+3   4.100225E+3   6.801171E-1   0.000000E+0   9.790571E-4   0.000000E+0   
9.865050E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.300286E+3   4.300286E+3   6.957529E-1   0.000000E+0   1.009175E-3   0.000000E+0   
9.990070E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.500161E+3   4.500161E+3   7.135960E-1   0.000000E+0   1.041487E-3   0.000000E+0   
1.011509E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.699982E+3   4.699982E+3   7.307067E-1   0.000000E+0   1.073062E-3   0.000000E+0   
1.024013E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.900140E+3   4.900140E+3   7.446276E-1   0.000000E+0   1.101472E-3   0.000000E+0   
1.036516E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.100248E+3   5.100248E+3   7.589922E-1   0.000000E+0   1.130322E-3   0.000000E+0   
1.049069E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.300048E+3   5.300048E+3   7.731229E-1   0.000000E+0   1.158916E-3   0.000000E+0   
1.061573E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.500009E+3   5.500009E+3   7.888226E-1   0.000000E+0   1.189090E-3   0.000000E+0   
1.074076E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.700173E+3   5.700173E+3   8.022165E-1   0.000000E+0   1.216974E-3   0.000000E+0   
1.086580E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.900313E+3   5.900313E+3   8.169553E-1   0.000000E+0   1.246200E-3   0.000000E+0   
1.099084E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.099977E+3   6.099977E+3   8.324042E-1   0.000000E+0   1.276103E-3   0.000000E+0   
1.111587E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.300217E+3   6.300217E+3   8.448552E-1   0.000000E+0   1.303049E-3   0.000000E+0   
1.124087E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.500296E+3   6.500296E+3   8.586595E-1   0.000000E+0   1.331336E-3   0.000000E+0   
1.136636E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.700114E+3   6.700114E+3   8.706756E-1   0.000000E+0   1.357817E-3   0.000000E+0   
1.149139E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.900139E+3   6.900139E+3   8.845961E-1   0.000000E+0   1.386217E-3   0.000000E+0   
1.161641E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.100315E+3   7.100315E+3   8.981087E-1   0.000000E+0   1.414220E-3   0.000000E+0   
1.174140E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.300280E+3   7.300280E+3   9.094652E-1   0.000000E+0   1.440051E-3   0.000000E+0   
1.186642E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.500208E+3   7.500208E+3   9.227839E-1   0.000000E+0   1.467843E-3   0.000000E+0   
1.199194E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.700105E+3   7.700105E+3   9.338533E-1   0.000000E+0   1.493382E-3   0.000000E+0   
1.211696E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.900037E+3   7.900037E+3   9.468394E-1   0.000000E+0   1.520841E-3   0.000000E+0   
1.224201E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.100170E+3   8.100170E+3   9.581633E-1   0.000000E+0   1.546652E-3   0.000000E+0   
1.236702E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.300349E+3   8.300349E+3   9.695974E-1   0.000000E+0   1.572577E-3   0.000000E+0   
1.249204E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.500224E+3   8.500224E+3   9.810776E-1   0.000000E+0   1.598526E-3   0.000000E+0   
1.261757E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.700246E+3   8.700246E+3   9.910582E-1   0.000000E+0   1.622986E-3   0.000000E+0   
1.274258E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.900235E+3   8.900235E+3   1.003389E+0   0.000000E+0   1.649793E-3   0.000000E+0   
1.286762E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.100361E+3   9.100361E+3   1.015117E+0   0.000000E+0   1.676008E-3   0.000000E+0   
1.299264E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.300308E+3   9.300308E+3   1.023568E+0   0.000000E+0   1.698932E-3   0.000000E+0   
1.311764E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.500079E+3   9.500079E+3   1.034775E+0   0.000000E+0   1.724601E-3   0.000000E+0   
1.324266E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.700019E+3   9.700019E+3   1.045734E+0   0.000000E+0   1.750033E-3   0.000000E+0   
1.336820E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.900173E+3   9.900173E+3   1.054645E+0   0.000000E+0   1.773433E-3   0.000000E+0   
1.349170E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000018E+4   1.000018E+4   1.059354E+0   0.000000E+0   1.785381E-3   0.000000E+0   
1.367613E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.199984E+4   1.199984E+4   1.148483E+0   0.000000E+0   2.019262E-3   0.000000E+0   
1.382314E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.399993E+4   1.399993E+4   1.221747E+0   0.000000E+0   2.237309E-3   0.000000E+0   
1.397017E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.599956E+4   1.599956E+4   1.279590E+0   0.000000E+0   2.440083E-3   0.000000E+0   
1.411720E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.799952E+4   1.799952E+4   1.328295E+0   0.000000E+0   2.633606E-3   0.000000E+0   
1.429711E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.599976E+4   1.599976E+4   1.283586E+0   0.000000E+0   2.444099E-3   0.000000E+0   
1.444415E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400025E+4   1.400025E+4   1.233510E+0   0.000000E+0   2.249096E-3   0.000000E+0   
1.459570E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200021E+4   1.200021E+4   1.180535E+0   0.000000E+0   2.051341E-3   0.000000E+0   
1.477570E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000013E+4   1.000013E+4   1.121594E+0   0.000000E+0   1.847618E-3   0.000000E+0   
1.493364E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.800326E+3   9.800326E+3   1.115241E+0   0.000000E+0   1.826801E-3   0.000000E+0   
1.505917E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.600376E+3   9.600376E+3   1.107606E+0   0.000000E+0   1.804692E-3   0.000000E+0   
1.518421E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.400082E+3   9.400082E+3   1.100558E+0   0.000000E+0   1.783145E-3   0.000000E+0   
1.530922E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.200193E+3   9.200193E+3   1.093784E+0   0.000000E+0   1.761902E-3   0.000000E+0   
1.543428E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.000386E+3   9.000386E+3   1.089263E+0   0.000000E+0   1.742917E-3   0.000000E+0   
1.555932E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.800064E+3   8.800064E+3   1.081329E+0   0.000000E+0   1.720482E-3   0.000000E+0   
1.568435E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.600242E+3   8.600242E+3   1.075610E+0   0.000000E+0   1.700298E-3   0.000000E+0   
1.580990E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.400135E+3   8.400135E+3   1.069322E+0   0.000000E+0   1.679525E-3   0.000000E+0   
1.593495E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.200284E+3   8.200284E+3   1.063312E+0   0.000000E+0   1.659048E-3   0.000000E+0   
1.605997E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.000331E+3   8.000331E+3   1.055428E+0   0.000000E+0   1.636690E-3   0.000000E+0   
1.618500E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.800212E+3   7.800212E+3   1.049118E+0   0.000000E+0   1.615893E-3   0.000000E+0   
1.631005E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.600062E+3   7.600062E+3   1.041890E+0   0.000000E+0   1.594177E-3   0.000000E+0   
1.643506E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.400215E+3   7.400215E+3   1.035027E+0   0.000000E+0   1.572847E-3   0.000000E+0   
1.656059E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.200233E+3   7.200233E+3   1.027161E+0   0.000000E+0   1.550505E-3   0.000000E+0   
1.668564E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.000168E+3   7.000168E+3   1.020985E+0   0.000000E+0   1.529846E-3   0.000000E+0   
1.681068E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.800075E+3   6.800075E+3   1.012892E+0   0.000000E+0   1.507269E-3   0.000000E+0   
1.693572E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.600082E+3   6.600082E+3   1.006514E+0   0.000000E+0   1.486414E-3   0.000000E+0   
1.706074E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.400167E+3   6.400167E+3   9.987720E-1   0.000000E+0   1.464201E-3   0.000000E+0   
1.718579E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.200185E+3   6.200185E+3   9.903178E-1   0.000000E+0   1.441270E-3   0.000000E+0   
1.731083E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.000317E+3   6.000317E+3   9.838374E-1   0.000000E+0   1.420322E-3   0.000000E+0   
1.743588E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.800242E+3   5.800242E+3   9.778883E-1   0.000000E+0   1.399889E-3   0.000000E+0   
1.756093E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.600016E+3   5.600016E+3   9.687933E-1   0.000000E+0   1.376300E-3   0.000000E+0   
1.768597E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.400091E+3   5.400091E+3   9.613273E-1   0.000000E+0   1.354362E-3   0.000000E+0   
1.781150E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.199947E+3   5.199947E+3   9.504217E-1   0.000000E+0   1.328969E-3   0.000000E+0   
1.793653E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.000047E+3   5.000047E+3   9.429166E-1   0.000000E+0   1.306993E-3   0.000000E+0   
1.806156E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.800154E+3   4.800154E+3   9.312102E-1   0.000000E+0   1.280817E-3   0.000000E+0   
1.818660E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.600200E+3   4.600200E+3   9.237267E-1   0.000000E+0   1.258859E-3   0.000000E+0   
1.831163E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.400186E+3   4.400186E+3   9.151202E-1   0.000000E+0   1.235774E-3   0.000000E+0   
1.843667E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.200250E+3   4.200250E+3   9.046928E-1   0.000000E+0   1.210873E-3   0.000000E+0   
1.856171E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.000182E+3   4.000182E+3   8.947223E-1   0.000000E+0   1.186420E-3   0.000000E+0   
1.868676E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.800035E+3   3.800035E+3   8.829697E-1   0.000000E+0   1.160179E-3   0.000000E+0   
1.881179E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.599884E+3   3.599884E+3   8.722821E-1   0.000000E+0   1.135003E-3   0.000000E+0   
1.893684E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.400013E+3   3.400013E+3   8.604485E-1   0.000000E+0   1.108701E-3   0.000000E+0   
1.906191E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.200195E+3   3.200195E+3   8.485079E-1   0.000000E+0   1.082296E-3   0.000000E+0   
1.918693E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.000191E+3   3.000191E+3   8.359051E-1   0.000000E+0   1.055216E-3   0.000000E+0   
1.931198E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.800065E+3   2.800065E+3   8.203858E-1   0.000000E+0   1.025210E-3   0.000000E+0   
1.943700E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.600201E+3   2.600201E+3   8.046605E-1   0.000000E+0   9.950164E-4   0.000000E+0   
1.956203E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.400161E+3   2.400161E+3   7.875827E-1   0.000000E+0   9.634580E-4   0.000000E+0   
1.968756E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.199832E+3   2.199832E+3   7.698908E-1   0.000000E+0   9.312646E-4   0.000000E+0   
1.981258E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.999885E+3   1.999885E+3   7.494180E-1   0.000000E+0   8.963181E-4   0.000000E+0   
1.993611E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.799974E+3   1.799974E+3   7.263983E-1   0.000000E+0   8.588272E-4   0.000000E+0   
2.005611E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.600146E+3   1.600146E+3   7.014615E-1   0.000000E+0   8.194252E-4   0.000000E+0   
2.017614E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400078E+3   1.400078E+3   6.721266E-1   0.000000E+0   7.756076E-4   0.000000E+0   
2.030067E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200067E+3   1.200067E+3   6.369890E-1   0.000000E+0   7.259915E-4   0.000000E+0   
2.042518E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.999160E+2   9.999160E+2   5.989169E-1   0.000000E+0   6.734310E-4   0.000000E+0   
2.054971E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.999372E+2   7.999372E+2   5.566816E-1   0.000000E+0   6.167195E-4   0.000000E+0   
2.067423E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.999011E+2   5.999011E+2   5.042527E-1   0.000000E+0   5.498103E-4   0.000000E+0   
2.079782E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.000083E+2   5.000083E+2   4.772924E-1   0.000000E+0   5.156190E-4   0.000000E+0   
2.095423E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.999616E+2   3.999616E+2   4.440854E-1   0.000000E+0   4.751698E-4   0.000000E+0   
2.107376E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.998077E+2   2.998077E+2   4.084424E-1   0.000000E+0   4.322768E-4   0.000000E+0   
2.119733E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.998469E+2   1.998469E+2   3.668522E-1   0.000000E+0   3.834506E-4   0.000000E+0   
2.131683E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000041E+2   1.000041E+2   3.194049E-1   0.000000E+0   3.287759E-4   0.000000E+0   
2.143483E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.391275E-1   -1.391275E-1   2.583518E-1   0.000000E+0   2.604736E-4   0.000000E+0   
2.155238E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.001107E+2   -1.001107E+2   1.869126E-1   0.000000E+0   1.817977E-4   0.000000E+0   
2.167040E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.001287E+2   -2.001287E+2   1.155593E-1   0.000000E+0   1.032042E-4   0.000000E+0   
2.178843E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.001038E+2   -3.001038E+2   5.292884E-2   0.000000E+0   3.333674E-5   0.000000E+0   
2.190644E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.000289E+2   -4.000289E+2   -5.031394E-3   0.000000E+0   -3.185690E-5   0.000000E+0   
2.202447E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.000683E+2   -5.000683E+2   -5.274810E-2   0.000000E+0   -8.681529E-5   0.000000E+0   
2.217585E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.000472E+2   -7.000472E+2   -1.350647E-1   0.000000E+0   -1.836080E-4   0.000000E+0   
2.229388E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.000511E+2   -9.000511E+2   -2.003095E-1   0.000000E+0   -2.633307E-4   0.000000E+0   
2.241191E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.100148E+3   -1.100148E+3   -2.518145E-1   0.000000E+0   -3.293204E-4   0.000000E+0   
2.253097E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.300170E+3   -1.300170E+3   -2.942410E-1   0.000000E+0   -3.862262E-4   0.000000E+0   
2.264998E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.500163E+3   -1.500163E+3   -3.317672E-1   0.000000E+0   -4.382295E-4   0.000000E+0   
2.276898E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.700224E+3   -1.700224E+3   -3.675856E-1   0.000000E+0   -4.885300E-4   0.000000E+0   
2.288800E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.900206E+3   -1.900206E+3   -3.998041E-1   0.000000E+0   -5.352248E-4   0.000000E+0   
2.300799E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.100157E+3   -2.100157E+3   -4.278912E-1   0.000000E+0   -5.777859E-4   0.000000E+0   
2.312752E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.300286E+3   -2.300286E+3   -4.555015E-1   0.000000E+0   -6.198833E-4   0.000000E+0   
2.324700E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.500093E+3   -2.500093E+3   -4.789292E-1   0.000000E+0   -6.577747E-4   0.000000E+0   
2.336599E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.700154E+3   -2.700154E+3   -4.999972E-1   0.000000E+0   -6.933248E-4   0.000000E+0   
2.348550E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.899993E+3   -2.899993E+3   -5.204346E-1   0.000000E+0   -7.282281E-4   0.000000E+0   
2.360496E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.100172E+3   -3.100172E+3   -5.427710E-1   0.000000E+0   -7.650551E-4   0.000000E+0   
2.372394E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.300101E+3   -3.300101E+3   -5.607776E-1   0.000000E+0   -7.975342E-4   0.000000E+0   
2.384345E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.500162E+3   -3.500162E+3   -5.832523E-1   0.000000E+0   -8.344910E-4   0.000000E+0   
2.396296E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.700012E+3   -3.700012E+3   -6.003697E-1   0.000000E+0   -8.660752E-4   0.000000E+0   
2.408245E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.900292E+3   -3.900292E+3   -6.198465E-1   0.000000E+0   -9.000498E-4   0.000000E+0   
2.420196E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.100160E+3   -4.100160E+3   -6.335231E-1   0.000000E+0   -9.281945E-4   0.000000E+0   
2.432147E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.300110E+3   -4.300110E+3   -6.521645E-1   0.000000E+0   -9.613100E-4   0.000000E+0   
2.444099E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.500167E+3   -4.500167E+3   -6.698444E-1   0.000000E+0   -9.934717E-4   0.000000E+0   
2.456049E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.700118E+3   -4.700118E+3   -6.844786E-1   0.000000E+0   -1.022580E-3   0.000000E+0   
2.467950E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.900089E+3   -4.900089E+3   -6.995370E-1   0.000000E+0   -1.052114E-3   0.000000E+0   
2.479899E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.100218E+3   -5.100218E+3   -7.157788E-1   0.000000E+0   -1.082843E-3   0.000000E+0   
2.491850E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.300151E+3   -5.300151E+3   -7.326122E-1   0.000000E+0   -1.114149E-3   0.000000E+0   
2.503802E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.500147E+3   -5.500147E+3   -7.450927E-1   0.000000E+0   -1.141107E-3   0.000000E+0   
2.515754E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.700298E+3   -5.700298E+3   -7.595874E-1   0.000000E+0   -1.170090E-3   0.000000E+0   
2.527705E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.900144E+3   -5.900144E+3   -7.733595E-1   0.000000E+0   -1.198329E-3   0.000000E+0   
2.539657E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.100145E+3   -6.100145E+3   -7.891484E-1   0.000000E+0   -1.228595E-3   0.000000E+0   
2.551604E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.300134E+3   -6.300134E+3   -7.995299E-1   0.000000E+0   -1.253454E-3   0.000000E+0   
2.563556E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.500024E+3   -6.500024E+3   -8.173491E-1   0.000000E+0   -1.285742E-3   0.000000E+0   
2.575506E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.700189E+3   -6.700189E+3   -8.285741E-1   0.000000E+0   -1.311457E-3   0.000000E+0   
2.587455E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.900253E+3   -6.900253E+3   -8.422330E-1   0.000000E+0   -1.339598E-3   0.000000E+0   
2.599356E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.100161E+3   -7.100161E+3   -8.521003E-1   0.000000E+0   -1.363937E-3   0.000000E+0   
2.611307E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.300275E+3   -7.300275E+3   -8.664619E-1   0.000000E+0   -1.392784E-3   0.000000E+0   
2.623256E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.500125E+3   -7.500125E+3   -8.802620E-1   0.000000E+0   -1.421051E-3   0.000000E+0   
2.635205E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.700022E+3   -7.700022E+3   -8.939670E-1   0.000000E+0   -1.449226E-3   0.000000E+0   
2.647105E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.900147E+3   -7.900147E+3   -9.035769E-1   0.000000E+0   -1.473323E-3   0.000000E+0   
2.659054E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.100094E+3   -8.100094E+3   -9.157333E-1   0.000000E+0   -1.499953E-3   0.000000E+0   
2.671007E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.300266E+3   -8.300266E+3   -9.266427E-1   0.000000E+0   -1.525352E-3   0.000000E+0   
2.682907E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.500263E+3   -8.500263E+3   -9.395471E-1   0.000000E+0   -1.552734E-3   0.000000E+0   
2.694857E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.700034E+3   -8.700034E+3   -9.514067E-1   0.000000E+0   -1.579055E-3   0.000000E+0   
2.706809E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.900228E+3   -8.900228E+3   -9.623549E-1   0.000000E+0   -1.604495E-3   0.000000E+0   
2.718753E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.100189E+3   -9.100189E+3   -9.719035E-1   0.000000E+0   -1.628518E-3   0.000000E+0   
2.730702E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.300200E+3   -9.300200E+3   -9.836639E-1   0.000000E+0   -1.654757E-3   0.000000E+0   
2.742708E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.500178E+3   -9.500178E+3   -9.954803E-1   0.000000E+0   -1.681050E-3   0.000000E+0   
2.754656E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.700107E+3   -9.700107E+3   -1.005061E+0   0.000000E+0   -1.705103E-3   0.000000E+0   
2.766607E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.900029E+3   -9.900029E+3   -1.015086E+0   0.000000E+0   -1.729600E-3   0.000000E+0   
2.778456E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.000012E+4   -1.000012E+4   -1.022097E+0   0.000000E+0   -1.743856E-3   0.000000E+0   
2.798007E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.199995E+4   -1.199995E+4   -1.115765E+0   0.000000E+0   -1.982289E-3   0.000000E+0   
2.812608E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.399974E+4   -1.399974E+4   -1.200430E+0   0.000000E+0   -2.211715E-3   0.000000E+0   
@@END Data.
@Time at end of measurement: 09:49:54
@NO Instrument  Changes.
@@Final Manipulated Data
New Section: Section 0: 
1.453500E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.399982E+4   -1.399982E+4   -1.161182E+0   0.000000E+0   5.220302E-4   0.000000E+0   
2.907600E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.199999E+4   -1.199999E+4   -1.106947E+0   0.000000E+0   3.361290E-4   0.000000E+0   
4.646500E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.000024E+4   -1.000024E+4   -1.059563E+0   0.000000E+0   1.433851E-4   0.000000E+0   
6.173500E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.800147E+3   -9.800147E+3   -1.048243E+0   0.000000E+0   1.306785E-4   0.000000E+0   
7.372300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.600204E+3   -9.600204E+3   -1.039898E+0   0.000000E+0   1.150140E-4   0.000000E+0   
8.566300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.400146E+3   -9.400146E+3   -1.034825E+0   0.000000E+0   9.606482E-5   0.000000E+0   
9.759500E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.200167E+3   -9.200167E+3   -1.030623E+0   0.000000E+0   7.625387E-5   0.000000E+0   
1.094890E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.000099E+3   -9.000099E+3   -1.024911E+0   0.000000E+0   5.794163E-5   0.000000E+0   
1.213770E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.800020E+3   -8.800020E+3   -1.020124E+0   0.000000E+0   3.870360E-5   0.000000E+0   
1.333700E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.600163E+3   -8.600163E+3   -1.014132E+0   0.000000E+0   2.069670E-5   0.000000E+0   
1.453090E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.400180E+3   -8.400180E+3   -1.008934E+0   0.000000E+0   1.880768E-6   0.000000E+0   
1.572460E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.200187E+3   -8.200187E+3   -1.000526E+0   0.000000E+0   -1.372621E-5   0.000000E+0   
1.691350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.000187E+3   -8.000187E+3   -9.954341E-1   0.000000E+0   -3.264986E-5   0.000000E+0   
1.810760E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.800201E+3   -7.800201E+3   -9.859596E-1   0.000000E+0   -4.718939E-5   0.000000E+0   
1.929640E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.600193E+3   -7.600193E+3   -9.827071E-1   0.000000E+0   -6.795357E-5   0.000000E+0   
2.049530E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.400190E+3   -7.400190E+3   -9.745225E-1   0.000000E+0   -8.378516E-5   0.000000E+0   
2.168960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.200254E+3   -7.200254E+3   -9.697457E-1   0.000000E+0   -1.030165E-4   0.000000E+0   
2.288350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.000128E+3   -7.000128E+3   -9.621676E-1   0.000000E+0   -1.194691E-4   0.000000E+0   
2.407780E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.800085E+3   -6.800085E+3   -9.558074E-1   0.000000E+0   -1.371299E-4   0.000000E+0   
2.527790E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.600138E+3   -6.600138E+3   -9.479659E-1   0.000000E+0   -1.532978E-4   0.000000E+0   
2.647310E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.400242E+3   -6.400242E+3   -9.418150E-1   0.000000E+0   -1.711502E-4   0.000000E+0   
2.766830E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.200156E+3   -6.200156E+3   -9.365604E-1   0.000000E+0   -1.899217E-4   0.000000E+0   
2.886350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.999998E+3   -5.999998E+3   -9.263450E-1   0.000000E+0   -2.037409E-4   0.000000E+0   
3.005840E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.800137E+3   -5.800137E+3   -9.211299E-1   0.000000E+0   -2.225249E-4   0.000000E+0   
3.125350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.600137E+3   -5.600137E+3   -9.105529E-1   0.000000E+0   -2.359636E-4   0.000000E+0   
3.244820E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.400026E+3   -5.400026E+3   -9.039486E-1   0.000000E+0   -2.533885E-4   0.000000E+0   
3.363850E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.200029E+3   -5.200029E+3   -8.969259E-1   0.000000E+0   -2.703811E-4   0.000000E+0   
3.483340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.000122E+3   -5.000122E+3   -8.889644E-1   0.000000E+0   -2.864242E-4   0.000000E+0   
3.602830E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.800043E+3   -4.800043E+3   -8.807722E-1   0.000000E+0   -3.022572E-4   0.000000E+0   
3.722340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.599999E+3   -4.599999E+3   -8.717974E-1   0.000000E+0   -3.173034E-4   0.000000E+0   
3.841340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.400078E+3   -4.400078E+3   -8.616852E-1   0.000000E+0   -3.311975E-4   0.000000E+0   
3.960860E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.199920E+3   -4.199920E+3   -8.523383E-1   0.000000E+0   -3.458853E-4   0.000000E+0   
4.080380E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.000027E+3   -4.000027E+3   -8.426935E-1   0.000000E+0   -3.602434E-4   0.000000E+0   
4.199910E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.800102E+3   -3.800102E+3   -8.317027E-1   0.000000E+0   -3.732594E-4   0.000000E+0   
4.319390E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.600044E+3   -3.600044E+3   -8.243541E-1   0.000000E+0   -3.899334E-4   0.000000E+0   
4.438910E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.399865E+3   -3.399865E+3   -8.096039E-1   0.000000E+0   -3.992205E-4   0.000000E+0   
4.558440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.200037E+3   -3.200037E+3   -7.974500E-1   0.000000E+0   -4.110618E-4   0.000000E+0   
4.677950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.000054E+3   -3.000054E+3   -7.852967E-1   0.000000E+0   -4.229221E-4   0.000000E+0   
4.797470E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.799954E+3   -2.799954E+3   -7.726228E-1   0.000000E+0   -4.342760E-4   0.000000E+0   
4.916970E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.600107E+3   -2.600107E+3   -7.603814E-1   0.000000E+0   -4.460320E-4   0.000000E+0   
5.036490E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.399867E+3   -2.399867E+3   -7.407769E-1   0.000000E+0   -4.504719E-4   0.000000E+0   
5.156000E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.199992E+3   -2.199992E+3   -7.228554E-1   0.000000E+0   -4.565512E-4   0.000000E+0   
5.276010E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.999931E+3   -1.999931E+3   -7.013866E-1   0.000000E+0   -4.591055E-4   0.000000E+0   
5.394020E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.799927E+3   -1.799927E+3   -6.802227E-1   0.000000E+0   -4.619578E-4   0.000000E+0   
5.513050E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.599884E+3   -1.599884E+3   -6.574467E-1   0.000000E+0   -4.632028E-4   0.000000E+0   
5.632050E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.400077E+3   -1.400077E+3   -6.274967E-1   0.000000E+0   -4.572454E-4   0.000000E+0   
5.751080E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.200030E+3   -1.200030E+3   -5.912459E-1   0.000000E+0   -4.450160E-4   0.000000E+0   
5.870090E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.998903E+2   -9.998903E+2   -5.564513E-1   0.000000E+0   -4.342538E-4   0.000000E+0   
5.988590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.999150E+2   -7.999150E+2   -5.104817E-1   0.000000E+0   -4.122970E-4   0.000000E+0   
6.107100E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.000578E+2   -6.000578E+2   -4.610431E-1   0.000000E+0   -3.868571E-4   0.000000E+0   
6.225100E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.998824E+2   -4.998824E+2   -4.297478E-1   0.000000E+0   -3.675907E-4   0.000000E+0   
6.375990E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.998894E+2   -3.998894E+2   -3.982557E-1   0.000000E+0   -3.481056E-4   0.000000E+0   
6.494010E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.998606E+2   -2.998606E+2   -3.632133E-1   0.000000E+0   -3.250745E-4   0.000000E+0   
6.612020E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.000107E+2   -2.000107E+2   -3.218639E-1   0.000000E+0   -2.957150E-4   0.000000E+0   
6.730040E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.992111E+1   -9.992111E+1   -2.736762E-1   0.000000E+0   -2.595459E-4   0.000000E+0   
6.848050E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.326898E-1   1.326898E-1   -2.119880E-1   0.000000E+0   -2.098720E-4   0.000000E+0   
6.971580E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.001579E+2   1.001579E+2   -1.397311E-1   0.000000E+0   -1.496261E-4   0.000000E+0   
7.095110E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.000328E+2   2.000328E+2   -7.114466E-2   0.000000E+0   -9.303247E-5   0.000000E+0   
7.215150E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.000866E+2   3.000866E+2   -7.578984E-3   0.000000E+0   -4.148113E-5   0.000000E+0   
7.338690E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.001655E+2   4.001655E+2   5.051231E-2   0.000000E+0   4.592821E-6   0.000000E+0   
7.458710E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.002193E+2   5.002193E+2   9.919279E-2   0.000000E+0   4.125897E-5   0.000000E+0   
7.615590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.002196E+2   7.002196E+2   1.791317E-1   0.000000E+0   9.718210E-5   0.000000E+0   
7.740120E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.000303E+2   9.000303E+2   2.448167E-1   0.000000E+0   1.388741E-4   0.000000E+0   
7.864650E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.100016E+3   1.100016E+3   2.979153E-1   0.000000E+0   1.679586E-4   0.000000E+0   
7.989180E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.300149E+3   1.300149E+3   3.398032E-1   0.000000E+0   1.858149E-4   0.000000E+0   
8.113710E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.499967E+3   1.499967E+3   3.793526E-1   0.000000E+0   2.013703E-4   0.000000E+0   
8.238240E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.700071E+3   1.700071E+3   4.138671E-1   0.000000E+0   2.118566E-4   0.000000E+0   
8.362840E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.900271E+3   1.900271E+3   4.454105E-1   0.000000E+0   2.193602E-4   0.000000E+0   
8.488360E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.100136E+3   2.100136E+3   4.743196E-1   0.000000E+0   2.242698E-4   0.000000E+0   
8.614380E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.300057E+3   2.300057E+3   4.980307E-1   0.000000E+0   2.239746E-4   0.000000E+0   
8.739400E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.500076E+3   2.500076E+3   5.208845E-1   0.000000E+0   2.228105E-4   0.000000E+0   
8.864450E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.700147E+3   2.700147E+3   5.482594E-1   0.000000E+0   2.261610E-4   0.000000E+0   
8.989500E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.900234E+3   2.900234E+3   5.692744E-1   0.000000E+0   2.231499E-4   0.000000E+0   
9.114530E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.100137E+3   3.100137E+3   5.869866E-1   0.000000E+0   2.168579E-4   0.000000E+0   
9.239580E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.299991E+3   3.299991E+3   6.064780E-1   0.000000E+0   2.123511E-4   0.000000E+0   
9.364590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.500299E+3   3.500299E+3   6.251796E-1   0.000000E+0   2.070000E-4   0.000000E+0   
9.489590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.700224E+3   3.700224E+3   6.443134E-1   0.000000E+0   2.021270E-4   0.000000E+0   
9.614560E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.900114E+3   3.900114E+3   6.607739E-1   0.000000E+0   1.945851E-4   0.000000E+0   
9.740040E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.100225E+3   4.100225E+3   6.801171E-1   0.000000E+0   1.898992E-4   0.000000E+0   
9.865050E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.300286E+3   4.300286E+3   6.957529E-1   0.000000E+0   1.815119E-4   0.000000E+0   
9.990070E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.500161E+3   4.500161E+3   7.135960E-1   0.000000E+0   1.753542E-4   0.000000E+0   
1.011509E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.699982E+3   4.699982E+3   7.307067E-1   0.000000E+0   1.684706E-4   0.000000E+0   
1.024013E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.900140E+3   4.900140E+3   7.446276E-1   0.000000E+0   1.583568E-4   0.000000E+0   
1.036516E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.100248E+3   5.100248E+3   7.589922E-1   0.000000E+0   1.486928E-4   0.000000E+0   
1.049069E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.300048E+3   5.300048E+3   7.731229E-1   0.000000E+0   1.388317E-4   0.000000E+0   
1.061573E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.500009E+3   5.500009E+3   7.888226E-1   0.000000E+0   1.305203E-4   0.000000E+0   
1.074076E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.700173E+3   5.700173E+3   8.022165E-1   0.000000E+0   1.198787E-4   0.000000E+0   
1.086580E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.900313E+3   5.900313E+3   8.169553E-1   0.000000E+0   1.105850E-4   0.000000E+0   
1.099084E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.099977E+3   6.099977E+3   8.324042E-1   0.000000E+0   1.020585E-4   0.000000E+0   
1.111587E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.300217E+3   6.300217E+3   8.448552E-1   0.000000E+0   9.046496E-5   0.000000E+0   
1.124087E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.500296E+3   6.500296E+3   8.586595E-1   0.000000E+0   8.024398E-5   0.000000E+0   
1.136636E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.700114E+3   6.700114E+3   8.706756E-1   0.000000E+0   6.826623E-5   0.000000E+0   
1.149139E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.900139E+3   6.900139E+3   8.845961E-1   0.000000E+0   5.816791E-5   0.000000E+0   
1.161641E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.100315E+3   7.100315E+3   8.981087E-1   0.000000E+0   4.764372E-5   0.000000E+0   
1.174140E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.300280E+3   7.300280E+3   9.094652E-1   0.000000E+0   3.498866E-5   0.000000E+0   
1.186642E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.500208E+3   7.500208E+3   9.227839E-1   0.000000E+0   2.430026E-5   0.000000E+0   
1.199194E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.700105E+3   7.700105E+3   9.338533E-1   0.000000E+0   1.136631E-5   0.000000E+0   
1.211696E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.900037E+3   7.900037E+3   9.468394E-1   0.000000E+0   3.447807E-7   0.000000E+0   
1.224201E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.100170E+3   8.100170E+3   9.581633E-1   0.000000E+0   -1.236299E-5   0.000000E+0   
1.236702E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.300349E+3   8.300349E+3   9.695974E-1   0.000000E+0   -2.496620E-5   0.000000E+0   
1.249204E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.500224E+3   8.500224E+3   9.810776E-1   0.000000E+0   -3.748669E-5   0.000000E+0   
1.261757E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.700246E+3   8.700246E+3   9.910582E-1   0.000000E+0   -5.152451E-5   0.000000E+0   
1.274258E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.900235E+3   8.900235E+3   1.003389E+0   0.000000E+0   -6.320843E-5   0.000000E+0   
1.286762E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.100361E+3   9.100361E+3   1.015117E+0   0.000000E+0   -7.551055E-5   0.000000E+0   
1.299264E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.300308E+3   9.300308E+3   1.023568E+0   0.000000E+0   -9.106971E-5   0.000000E+0   
1.311764E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.500079E+3   9.500079E+3   1.034775E+0   0.000000E+0   -1.038505E-4   0.000000E+0   
1.324266E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.700019E+3   9.700019E+3   1.045734E+0   0.000000E+0   -1.169001E-4   0.000000E+0   
1.336820E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.900173E+3   9.900173E+3   1.054645E+0   0.000000E+0   -1.320231E-4   0.000000E+0   
1.349170E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000018E+4   1.000018E+4   1.059354E+0   0.000000E+0   -1.393230E-4   0.000000E+0   
1.367613E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.199984E+4   1.199984E+4   1.148483E+0   0.000000E+0   -2.903111E-4   0.000000E+0   
1.382314E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.399993E+4   1.399993E+4   1.221747E+0   0.000000E+0   -4.572156E-4   0.000000E+0   
1.397017E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.599956E+4   1.599956E+4   1.279590E+0   0.000000E+0   -6.347811E-4   0.000000E+0   
1.411720E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.799952E+4   1.799952E+4   1.328295E+0   0.000000E+0   -8.078257E-4   0.000000E+0   
1.429711E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.599976E+4   1.599976E+4   1.283586E+0   0.000000E+0   -6.308014E-4   0.000000E+0   
1.444415E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400025E+4   1.400025E+4   1.233510E+0   0.000000E+0   -4.454903E-4   0.000000E+0   
1.459570E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200021E+4   1.200021E+4   1.180535E+0   0.000000E+0   -2.583034E-4   0.000000E+0   
1.477570E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000013E+4   1.000013E+4   1.121594E+0   0.000000E+0   -7.707631E-5   0.000000E+0   
1.493364E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.800326E+3   9.800326E+3   1.115241E+0   0.000000E+0   -5.943790E-5   0.000000E+0   
1.505917E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.600376E+3   9.600376E+3   1.107606E+0   0.000000E+0   -4.306357E-5   0.000000E+0   
1.518421E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.400082E+3   9.400082E+3   1.100558E+0   0.000000E+0   -2.606040E-5   0.000000E+0   
1.530922E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.200193E+3   9.200193E+3   1.093784E+0   0.000000E+0   -8.831846E-6   0.000000E+0   
1.543428E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.000386E+3   9.000386E+3   1.089263E+0   0.000000E+0   1.063948E-5   0.000000E+0   
1.555932E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.800064E+3   8.800064E+3   1.081329E+0   0.000000E+0   2.676058E-5   0.000000E+0   
1.568435E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.600242E+3   8.600242E+3   1.075610E+0   0.000000E+0   4.503559E-5   0.000000E+0   
1.580990E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.400135E+3   8.400135E+3   1.069322E+0   0.000000E+0   6.277599E-5   0.000000E+0   
1.593495E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.200284E+3   8.200284E+3   1.063312E+0   0.000000E+0   8.076358E-5   0.000000E+0   
1.605997E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.000331E+3   8.000331E+3   1.055428E+0   0.000000E+0   9.689047E-5   0.000000E+0   
1.618500E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.800212E+3   7.800212E+3   1.049118E+0   0.000000E+0   1.146097E-4   0.000000E+0   
1.631005E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.600062E+3   7.600062E+3   1.041890E+0   0.000000E+0   1.314156E-4   0.000000E+0   
1.643506E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.400215E+3   7.400215E+3   1.035027E+0   0.000000E+0   1.485499E-4   0.000000E+0   
1.656059E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.200233E+3   7.200233E+3   1.027161E+0   0.000000E+0   1.646976E-4   0.000000E+0   
1.668564E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.000168E+3   7.000168E+3   1.020985E+0   0.000000E+0   1.825451E-4   0.000000E+0   
1.681068E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.800075E+3   6.800075E+3   1.012892E+0   0.000000E+0   1.984793E-4   0.000000E+0   
1.693572E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.600082E+3   6.600082E+3   1.006514E+0   0.000000E+0   2.161163E-4   0.000000E+0   
1.706074E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.400167E+3   6.400167E+3   9.987720E-1   0.000000E+0   2.323798E-4   0.000000E+0   
1.718579E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.200185E+3   6.200185E+3   9.903178E-1   0.000000E+0   2.479393E-4   0.000000E+0   
1.731083E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.000317E+3   6.000317E+3   9.838374E-1   0.000000E+0   2.654588E-4   0.000000E+0   
1.743588E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.800242E+3   5.800242E+3   9.778883E-1   0.000000E+0   2.835345E-4   0.000000E+0   
1.756093E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.600016E+3   5.600016E+3   9.687933E-1   0.000000E+0   2.984823E-4   0.000000E+0   
1.768597E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.400091E+3   5.400091E+3   9.613273E-1   0.000000E+0   3.150231E-4   0.000000E+0   
1.781150E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.199947E+3   5.199947E+3   9.504217E-1   0.000000E+0   3.281505E-4   0.000000E+0   
1.793653E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.000047E+3   5.000047E+3   9.429166E-1   0.000000E+0   3.446491E-4   0.000000E+0   
1.806156E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.800154E+3   4.800154E+3   9.312102E-1   0.000000E+0   3.569456E-4   0.000000E+0   
1.818660E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.600200E+3   4.600200E+3   9.237267E-1   0.000000E+0   3.734723E-4   0.000000E+0   
1.831163E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.400186E+3   4.400186E+3   9.151202E-1   0.000000E+0   3.888833E-4   0.000000E+0   
1.843667E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.200250E+3   4.200250E+3   9.046928E-1   0.000000E+0   4.024640E-4   0.000000E+0   
1.856171E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.000182E+3   4.000182E+3   8.947223E-1   0.000000E+0   4.165174E-4   0.000000E+0   
1.868676E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.800035E+3   3.800035E+3   8.829697E-1   0.000000E+0   4.287982E-4   0.000000E+0   
1.881179E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.599884E+3   3.599884E+3   8.722821E-1   0.000000E+0   4.421444E-4   0.000000E+0   
1.893684E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.400013E+3   3.400013E+3   8.604485E-1   0.000000E+0   4.543112E-4   0.000000E+0   
1.906191E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.200195E+3   3.200195E+3   8.485079E-1   0.000000E+0   4.663645E-4   0.000000E+0   
1.918693E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.000191E+3   3.000191E+3   8.359051E-1   0.000000E+0   4.777779E-4   0.000000E+0   
1.931198E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.800065E+3   2.800065E+3   8.203858E-1   0.000000E+0   4.862894E-4   0.000000E+0   
1.943700E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.600201E+3   2.600201E+3   8.046605E-1   0.000000E+0   4.945635E-4   0.000000E+0   
1.956203E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.400161E+3   2.400161E+3   7.875827E-1   0.000000E+0   5.015062E-4   0.000000E+0   
1.968756E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.199832E+3   2.199832E+3   7.698908E-1   0.000000E+0   5.078696E-4   0.000000E+0   
1.981258E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.999885E+3   1.999885E+3   7.494180E-1   0.000000E+0   5.114062E-4   0.000000E+0   
1.993611E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.799974E+3   1.799974E+3   7.263983E-1   0.000000E+0   5.123915E-4   0.000000E+0   
2.005611E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.600146E+3   1.600146E+3   7.014615E-1   0.000000E+0   5.114499E-4   0.000000E+0   
2.017614E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400078E+3   1.400078E+3   6.721266E-1   0.000000E+0   5.061389E-4   0.000000E+0   
2.030067E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200067E+3   1.200067E+3   6.369890E-1   0.000000E+0   4.950184E-4   0.000000E+0   
2.042518E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.999160E+2   9.999160E+2   5.989169E-1   0.000000E+0   4.809802E-4   0.000000E+0   
2.054971E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.999372E+2   7.999372E+2   5.566816E-1   0.000000E+0   4.627580E-4   0.000000E+0   
2.067423E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.999011E+2   5.999011E+2   5.042527E-1   0.000000E+0   4.343492E-4   0.000000E+0   
2.079782E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.000083E+2   5.000083E+2   4.772924E-1   0.000000E+0   4.193839E-4   0.000000E+0   
2.095423E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.999616E+2   3.999616E+2   4.440854E-1   0.000000E+0   3.981904E-4   0.000000E+0   
2.107376E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.998077E+2   2.998077E+2   4.084424E-1   0.000000E+0   3.745737E-4   0.000000E+0   
2.119733E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.998469E+2   1.998469E+2   3.668522E-1   0.000000E+0   3.449867E-4   0.000000E+0   
2.131683E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000041E+2   1.000041E+2   3.194049E-1   0.000000E+0   3.095284E-4   0.000000E+0   
2.143483E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.391275E-1   -1.391275E-1   2.583518E-1   0.000000E+0   2.605004E-4   0.000000E+0   
2.155238E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.001107E+2   -1.001107E+2   1.869126E-1   0.000000E+0   2.010657E-4   0.000000E+0   
2.167040E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.001287E+2   -2.001287E+2   1.155593E-1   0.000000E+0   1.417224E-4   0.000000E+0   
2.178843E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.001038E+2   -3.001038E+2   5.292884E-2   0.000000E+0   9.109681E-5   0.000000E+0   
2.190644E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.000289E+2   -4.000289E+2   -5.031394E-3   0.000000E+0   4.513545E-5   0.000000E+0   
2.202447E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.000683E+2   -5.000683E+2   -5.274810E-2   0.000000E+0   9.431353E-6   0.000000E+0   
2.217585E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.000472E+2   -7.000472E+2   -1.350647E-1   0.000000E+0   -4.887201E-5   0.000000E+0   
2.229388E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.000511E+2   -9.000511E+2   -2.003095E-1   0.000000E+0   -9.010061E-5   0.000000E+0   
2.241191E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.100148E+3   -1.100148E+3   -2.518145E-1   0.000000E+0   -1.175783E-4   0.000000E+0   
2.253097E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.300170E+3   -1.300170E+3   -2.942410E-1   0.000000E+0   -1.359864E-4   0.000000E+0   
2.264998E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.500163E+3   -1.500163E+3   -3.317672E-1   0.000000E+0   -1.494977E-4   0.000000E+0   
2.276898E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.700224E+3   -1.700224E+3   -3.675856E-1   0.000000E+0   -1.612930E-4   0.000000E+0   
2.288800E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.900206E+3   -1.900206E+3   -3.998041E-1   0.000000E+0   -1.694978E-4   0.000000E+0   
2.300799E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.100157E+3   -2.100157E+3   -4.278912E-1   0.000000E+0   -1.735751E-4   0.000000E+0   
2.312752E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.300286E+3   -2.300286E+3   -4.555015E-1   0.000000E+0   -1.771542E-4   0.000000E+0   
2.324700E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.500093E+3   -2.500093E+3   -4.789292E-1   0.000000E+0   -1.765894E-4   0.000000E+0   
2.336599E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.700154E+3   -2.700154E+3   -4.999972E-1   0.000000E+0   -1.736343E-4   0.000000E+0   
2.348550E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.899993E+3   -2.899993E+3   -5.204346E-1   0.000000E+0   -1.700752E-4   0.000000E+0   
2.360496E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.100172E+3   -3.100172E+3   -5.427710E-1   0.000000E+0   -1.683743E-4   0.000000E+0   
2.372394E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.300101E+3   -3.300101E+3   -5.607776E-1   0.000000E+0   -1.623737E-4   0.000000E+0   
2.384345E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.500162E+3   -3.500162E+3   -5.832523E-1   0.000000E+0   -1.608253E-4   0.000000E+0   
2.396296E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.700012E+3   -3.700012E+3   -6.003697E-1   0.000000E+0   -1.539450E-4   0.000000E+0   
2.408245E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.900292E+3   -3.900292E+3   -6.198465E-1   0.000000E+0   -1.493725E-4   0.000000E+0   
2.420196E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.100160E+3   -4.100160E+3   -6.335231E-1   0.000000E+0   -1.390492E-4   0.000000E+0   
2.432147E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.300110E+3   -4.300110E+3   -6.521645E-1   0.000000E+0   -1.336809E-4   0.000000E+0   
2.444099E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.500167E+3   -4.500167E+3   -6.698444E-1   0.000000E+0   -1.273381E-4   0.000000E+0   
2.456049E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.700118E+3   -4.700118E+3   -6.844786E-1   0.000000E+0   -1.179626E-4   0.000000E+0   
2.467950E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.900089E+3   -4.900089E+3   -6.995370E-1   0.000000E+0   -1.090086E-4   0.000000E+0   
2.479899E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.100218E+3   -5.100218E+3   -7.157788E-1   0.000000E+0   -1.012191E-4   0.000000E+0   
2.491850E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.300151E+3   -5.300151E+3   -7.326122E-1   0.000000E+0   -9.404492E-5   0.000000E+0   
2.503802E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.500147E+3   -5.500147E+3   -7.450927E-1   0.000000E+0   -8.251003E-5   0.000000E+0   
2.515754E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.700298E+3   -5.700298E+3   -7.595874E-1   0.000000E+0   -7.297098E-5   0.000000E+0   
2.527705E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.900144E+3   -5.900144E+3   -7.733595E-1   0.000000E+0   -6.274576E-5   0.000000E+0   
2.539657E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.100145E+3   -6.100145E+3   -7.891484E-1   0.000000E+0   -5.451884E-5   0.000000E+0   
2.551604E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.300134E+3   -6.300134E+3   -7.995299E-1   0.000000E+0   -4.088587E-5   0.000000E+0   
2.563556E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.500024E+3   -6.500024E+3   -8.173491E-1   0.000000E+0   -3.470254E-5   0.000000E+0   
2.575506E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.700189E+3   -6.700189E+3   -8.285741E-1   0.000000E+0   -2.189199E-5   0.000000E+0   
2.587455E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.900253E+3   -6.900253E+3   -8.422330E-1   0.000000E+0   -1.152739E-5   0.000000E+0   
2.599356E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.100161E+3   -7.100161E+3   -8.521003E-1   0.000000E+0   2.609879E-6   0.000000E+0   
2.611307E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.300275E+3   -7.300275E+3   -8.664619E-1   0.000000E+0   1.227780E-5   0.000000E+0   
2.623256E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.500125E+3   -7.500125E+3   -8.802620E-1   0.000000E+0   2.247548E-5   0.000000E+0   
2.635205E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.700022E+3   -7.700022E+3   -8.939670E-1   0.000000E+0   3.277386E-5   0.000000E+0   
2.647105E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.900147E+3   -7.900147E+3   -9.035769E-1   0.000000E+0   4.719470E-5   0.000000E+0   
2.659054E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.100094E+3   -8.100094E+3   -9.157333E-1   0.000000E+0   5.904771E-5   0.000000E+0   
2.671007E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.300266E+3   -8.300266E+3   -9.266427E-1   0.000000E+0   7.217471E-5   0.000000E+0   
2.682907E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.500263E+3   -8.500263E+3   -9.395471E-1   0.000000E+0   8.328558E-5   0.000000E+0   
2.694857E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.700034E+3   -8.700034E+3   -9.514067E-1   0.000000E+0   9.541430E-5   0.000000E+0   
2.706809E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.900228E+3   -8.900228E+3   -9.623549E-1   0.000000E+0   1.085051E-4   0.000000E+0   
2.718753E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.100189E+3   -9.100189E+3   -9.719035E-1   0.000000E+0   1.229676E-4   0.000000E+0   
2.730702E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.300200E+3   -9.300200E+3   -9.836639E-1   0.000000E+0   1.352242E-4   0.000000E+0   
2.742708E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.500178E+3   -9.500178E+3   -9.954803E-1   0.000000E+0   1.474210E-4   0.000000E+0   
2.754656E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.700107E+3   -9.700107E+3   -1.005061E+0   0.000000E+0   1.618471E-4   0.000000E+0   
2.766607E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.900029E+3   -9.900029E+3   -1.015086E+0   0.000000E+0   1.758290E-4   0.000000E+0   
2.778456E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.000012E+4   -1.000012E+4   -1.022097E+0   0.000000E+0   1.808363E-4   0.000000E+0   
2.798007E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.199995E+4   -1.199995E+4   -1.115765E+0   0.000000E+0   3.273052E-4   0.000000E+0   
2.812608E+3   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.399974E+4   -1.399974E+4   -1.200430E+0   0.000000E+0   4.827723E-4   0.000000E+0   
@@END Data.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -13999.820     -13999.738     -0.041         Coercive Field: Field at which M//H changes sign
Ms emu                                  522.030E-6     -807.826E-6    664.928E-6     Saturation Magnetization: maximum M measured
Hc offset Oe                            -13999.82      -13999.74      -13999.78      (Hc upward curve + Hc Downward curve)/2 
M at H max emu                          -807.826E-6    522.030E-6     664.928E-6     M at the maximum field                  
PP emu                                  1.330E-3       1.143E-3       1.330E-3       Peak to Peak Signal (Max - Min)         
Stdev emu                               247.080E-6     242.456E-6     265.168E-6     Standard Deviation                      
Mr emu                                  -209.938E-6    260.568E-6     235.253E-6     Remanent Magnetization: M at H=0        
                                                                                                                             
HcP1                                    -17999.523     -17999.523     0.000          Pin 1 coercive field                    
HcP2                                    400.029        399.889        0.070          Pin 2 coercive field                    

@END Measurement parameters
